[aimspice]
[description]
3157
* This is a parametrized testbench for your pixel circuit array

* You should at least test your circuit with:
*	- current of 50 pA and exposure time 30 ms
*	- current of 750 pA and exposure time 2 ms

* Instructions
* Connect EXPOSE, ERASE, NRE_R1 and NRE_R2 at the right place
* Run a transient simulation with length 60 ms
* Make sure outputs of pixel circuits to ADC are called OUT1 and OUT2
* Make plots of output voltages to ADC (here called OUT1 and OUT2)
* The voltage across internal capacitor (any pixel) is also of interest (here called OUT_SAMPLED1)
* You should also plot the control signals EXPOSE, NRE_R1, NRE_R2 and ERASE

.include F:\AIMspice-simulations\Project\p18_cmos_models_tt.inc

* --------- Simulation Paramters ---------
.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(OUT1) V(OUT2) V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE) V(P11:N2)
.plot V(OUT_SAMPLED1)

* --------- Component Paramters ---------
.param LM124 = 1.08u
.param WM124 = 1.08u
.param LM3 = 1.08u
.param WM3 = 5.04u
.param LMC = 0.36u
.param WMC = 5.04u
.param C_CS = 2.5p
.param C_CC = 3p

* --------- Photodiode --------- 
.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1            ! Photo current source
d1 N1_R1C1 VDD dwell 1                        ! Reverse biased Diode
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40 ! Diode model
Cd1 N1_R1C1 VDD 30f                           ! Photo diode capacitor
.ends

* --------- Individual pixel circuit ---------
.subckt PixelCircuit VDD VSS OUT EXPOSE ERASE NRE
XPhoto VDD N1 PhotoDiode
M1 N1 EXPOSE N2 VSS NMOS L=LM124 W=WM124
M2 N2 ERASE VSS VSS NMOS L=LM124 W=WM124
CS N2 VSS C_CS
M3 VSS N2 N3 VDD PMOS L=LM3 W=WM3
M4 N3 NRE OUT VDD PMOS L=LM124 W=WM124
.ends

* --------- 4 pixel circuit ---------
MC1 OUT1 OUT1 1 1 PMOS L=LMC W=WMC
MC2 OUT2 OUT2 1 1 PMOS L=LMC W=WMC
CC1 OUT1 0 C_CC
CC2 OUT2 0 C_CC
XP11 1 0 OUT1 EXPOSE ERASE NRE_R1 PixelCircuit
XP12 1 0 OUT2 EXPOSE ERASE NRE_R1 PixelCircuit
XP21 1 0 OUT1 EXPOSE ERASE NRE_R2 PixelCircuit
XP22 1 0 OUT2 EXPOSE ERASE NRE_R2 PixelCircuit




[tran]
0.1ms
60ms
X
X
0
[ana]
4 0
[end]
