module FSM_ex_control (input wire Init, Clk, Reset